*** SPICE deck for cell Capacitance_Sim{sch} from library Project1
*** Created on Fri Jul 02, 2021 14:14:54
*** Last revised on Sat Jul 03, 2021 04:29:21
*** Written on Sat Jul 03, 2021 04:30:18 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: Capacitance_Sim{sch}
Mnmos@0 OUT net@9 gnd gnd NMOS L=0.14U W=0.21U
Mpmos@0 vdd net@9 OUT vdd PMOS L=0.14U W=0.49U
Rres@0 net@9 IN 20k

* Spice Code nodes in cell cell 'Capacitance_Sim{sch}'
vdd vdd gnd dc 1.8
vin In gnd (pulse 0 1.8 0.000001ns 0.000001ns 0.000001ns 10ns)
.tran 0.01ns 30.5ns
.include /home/nada/Desktop/DD2_Project1/130nm_bulk.pm
.control
run
set color0=white
set color1=black
set xbrushwidth=2
plot v(in) v(out)
.endc
.END
