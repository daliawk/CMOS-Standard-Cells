*** SPICE deck for cell NOR_1_Cinv_sim{sch} from library Project1
*** Created on Sun Jul 04, 2021 22:30:41
*** Last revised on Mon Jul 05, 2021 01:28:56
*** Written on Mon Jul 05, 2021 01:28:59 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Project1__INV_1 FROM CELL INV_1{sch}
.SUBCKT Project1__INV_1 gnd IN OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT IN gnd gnd NMOS L=0.14U W=0.21U
Mpmos@0 vdd IN OUT vdd PMOS L=0.14U W=0.49U
.ENDS Project1__INV_1

*** SUBCIRCUIT Project1__NOR_1 FROM CELL NOR_1{sch}
.SUBCKT Project1__NOR_1 gnd IN1 IN2 OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT IN2 gnd gnd nmos L=0.14U W=0.21U
Mnmos@1 OUT IN1 gnd gnd nmos' L=0.14U W=0.21U
Mpmos@0 vdd IN1 net@0 vdd pmos L=0.14U W=0.98U
Mpmos@1 net@0 IN2 OUT vdd pmos L=0.14U W=0.98U
.ENDS Project1__NOR_1

.global gnd vdd

*** TOP LEVEL CELL: NOR_1_Cinv_sim{sch}
XINV_1@0 gnd OUT INV_1@0_OUT vdd Project1__INV_1
XNOR_1@0 gnd IN1 IN2 OUT vdd Project1__NOR_1

* Spice Code nodes in cell cell 'NOR_1_Cinv_sim{sch}'
vdd VDD GND dc 1.8
vin1 IN1 gnd pulse(0 1.8 5000ps 0ps 0ps 5000ps)
vin2 IN2 gnd pulse(0 1.8 5000ps 0ps 0ps 5000ps)
.tran 10ns 50ns
.meas TRAN tpdf TRIG V(IN1) val=0.9 rise=1 TARG V(OUT) val=1.7 fall=1
.meas TRAN tpdr TRIG V(IN1) val=0.9 fall=1 TARG V(OUT) val=1.7 rise=1
.include /home/daliawk/DD2_Project1/130nm_bulk.pm
.control
run
set color0=white
set color1=black
set xbrushwidth=2
plot v(IN1) v(IN2) v(OUT)
.endc
.END
