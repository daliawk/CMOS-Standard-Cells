*** SPICE deck for cell INV_1_sim{sch} from library Project1
*** Created on Sat Jul 03, 2021 05:02:36
*** Last revised on Sat Jul 03, 2021 05:52:28
*** Written on Sat Jul 03, 2021 05:52:36 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Project1__INV_1 FROM CELL INV_1{sch}
.SUBCKT Project1__INV_1 gnd IN OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT IN gnd gnd NMOS L=0.14U W=0.21U
Mpmos@0 vdd IN OUT vdd PMOS L=0.14U W=0.49U
.ENDS Project1__INV_1

.global gnd vdd

*** TOP LEVEL CELL: INV_1_sim{sch}
Ccap@0 gnd OUT 2.17f
XINV_1@0 gnd INV_1@0_IN OUT vdd Project1__INV_1

* Spice Code nodes in cell cell 'INV_1_sim{sch}'
vdd VDD GND dc 1.8
vin IN gnd (pulse 0 1.8 500ps 480ps 480ps 1000ps)
.tran 10ps 3000ps
.meas TRAN tpdf TRIG V(IN) val=0.9 rise=1 TARG V(OUT) val=0.9 fall=1
.meas TRAN tpdr TRIG V(IN) val=0.9 fall=1 TARG V(OUT) val=0.9 rise=1
.include /home/nada/Desktop/DD2_Project1/130nm_bulk.pm
.control
run
set color0=white
set color1=black
set xbrushwidth=2
plot v(IN) v(OUT)
.endc
.END
