*** SPICE deck for cell COMPLEX_1_Cinv_Sim{sch} from library Project1
*** Created on Mon Jul 05, 2021 01:30:55
*** Last revised on Mon Jul 05, 2021 01:36:17
*** Written on Mon Jul 05, 2021 01:36:20 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Project1__COMPLEX_1 FROM CELL COMPLEX_1{sch}
.SUBCKT Project1__COMPLEX_1 gnd IN1 IN2 IN3 OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT IN1 net@16 gnd nmos L=0.14U W=0.42U
Mnmos@1 net@16 IN2 gnd gnd nmos L=0.14U W=0.42U
Mnmos@2 net@80 IN1 gnd gnd nmos L=0.14U W=0.42U
Mnmos@3 net@80 IN2 gnd gnd nmos L=0.14U W=0.42U
Mnmos@4 OUT IN3 net@80 gnd nmos L=0.14U W=0.42U
Mpmos@0 vdd IN2 net@0 vdd pmos L=0.14U W=0.98U
Mpmos@1 net@0 IN1 OUT vdd pmos L=0.14U W=0.98U
Mpmos@2 vdd IN1 net@10 vdd pmos L=0.14U W=0.98U
Mpmos@3 vdd IN2 net@10 vdd pmos L=0.14U W=0.98U
Mpmos@4 net@10 IN3 OUT vdd pmos L=0.14U W=0.98U
.ENDS Project1__COMPLEX_1

*** SUBCIRCUIT Project1__INV_1 FROM CELL INV_1{sch}
.SUBCKT Project1__INV_1 gnd IN OUT vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 OUT IN gnd gnd NMOS L=0.14U W=0.21U
Mpmos@0 vdd IN OUT vdd PMOS L=0.14U W=0.49U
.ENDS Project1__INV_1

.global gnd vdd

*** TOP LEVEL CELL: COMPLEX_1_Cinv_Sim{sch}
XCOMPLEX_@0 gnd IN1 IN2 IN3 OUT vdd Project1__COMPLEX_1
XINV_1@0 gnd OUT INV_1@0_OUT vdd Project1__INV_1

* Spice Code nodes in cell cell 'COMPLEX_1_Cinv_Sim{sch}'
vdd VDD GND dc 1.8
vin1 IN1 gnd pulse(0 1.8 5000ps 0ps 0ps 5000ps)
vin2 IN2 gnd pulse(0 1.8 5000ps 0ps 0ps 5000ps)
vin3 IN3 gnd pulse(0 0 5000ps 0ps 0ps 5000ps)
.tran 10ns 50ns
.meas TRAN tpdf TRIG V(IN1) val=0.9 rise=1 TARG V(OUT) val= 0.9 fall=1
.meas TRAN tpdr TRIG V(IN1) val=0.9 fall=1 TARG V(OUT) val=0.9 rise=1
.include /home/daliawk/DD2_Project1/130nm_bulk.pm
.control
run
set color0=white
set color1=black
set xbrushwidth=2
plot v(IN1) v(IN2) v(OUT)
.endc
.END
